// vga_char_params.vh
`ifndef VGA_CHAR_PARAMS_VH
`define VGA_CHAR_PARAMS_VH

//num_zero- num_nine: 32x32 pixel font for numbers 0-9

//char_dai:待
//char_ding:定
//char_mo:模
//char_shi:式
//char_ji:计
//char_suan:算
//char_xue:学
//char_xi:习
//char_yan:演
//char_shi2:示
//char_dui:对
//char_cuo:错

parameter num_zero={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11111000, 0b00000000, 0b00000000, 
    0b00001111, 0b11111110, 0b00000000, 0b00000000, 
    0b00001111, 0b11111111, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b00000000, 0b00000000, 
    0b00111110, 0b00001111, 0b10000000, 0b00000000, 
    0b00111100, 0b00000111, 0b10000000, 0b00000000, 
    0b00111100, 0b00000111, 0b11000000, 0b00000000, 
    0b01111100, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111100, 0b00000011, 0b11000000, 0b00000000, 
    0b00111100, 0b00000111, 0b10000000, 0b00000000, 
    0b00111110, 0b00000111, 0b10000000, 0b00000000, 
    0b00111111, 0b00001111, 0b10000000, 0b00000000, 
    0b00011111, 0b11111111, 0b00000000, 0b00000000, 
    0b00001111, 0b11111111, 0b00000000, 0b00000000, 
    0b00000111, 0b11111100, 0b00000000, 0b00000000, 
    0b00000001, 0b11111000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter num_one={
     0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000001, 0b11000000, 0b00000000, 0b00000000, 
    0b00000111, 0b11000000, 0b00000000, 0b00000000, 
    0b00001111, 0b11000000, 0b00000000, 0b00000000, 
    0b00111111, 0b11000000, 0b00000000, 0b00000000, 
    0b01111111, 0b11000000, 0b00000000, 0b00000000, 
    0b01111111, 0b11000000, 0b00000000, 0b00000000, 
    0b01111011, 0b11000000, 0b00000000, 0b00000000, 
    0b01100011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter num_two={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11111100, 0b00000000, 0b00000000, 
    0b00000111, 0b11111110, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b10000000, 0b00000000, 
    0b00111110, 0b00000111, 0b10000000, 0b00000000, 
    0b00111110, 0b00000111, 0b11000000, 0b00000000, 
    0b00111100, 0b00000011, 0b11000000, 0b00000000, 
    0b00111100, 0b00000011, 0b11000000, 0b00000000, 
    0b00111100, 0b00000111, 0b11000000, 0b00000000, 
    0b00111000, 0b00000111, 0b10000000, 0b00000000, 
    0b00000000, 0b00001111, 0b10000000, 0b00000000, 
    0b00000000, 0b00011111, 0b10000000, 0b00000000, 
    0b00000000, 0b00111111, 0b00000000, 0b00000000, 
    0b00000000, 0b11111110, 0b00000000, 0b00000000, 
    0b00000001, 0b11111100, 0b00000000, 0b00000000, 
    0b00000011, 0b11111000, 0b00000000, 0b00000000, 
    0b00000111, 0b11100000, 0b00000000, 0b00000000, 
    0b00001111, 0b11000000, 0b00000000, 0b00000000, 
    0b00011111, 0b10000000, 0b00000000, 0b00000000, 
    0b00111111, 0b00000000, 0b00000000, 0b00000000, 
    0b00111110, 0b00000000, 0b00000000, 0b00000000, 
    0b00111111, 0b11111111, 0b11000000, 0b00000000, 
    0b01111111, 0b11111111, 0b11000000, 0b00000000, 
    0b01111111, 0b11111111, 0b11000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter num_three={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11111100, 0b00000000, 0b00000000, 
    0b00001111, 0b11111111, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b10000000, 0b00000000, 
    0b00111110, 0b00000111, 0b10000000, 0b00000000, 
    0b00111100, 0b00000111, 0b11000000, 0b00000000, 
    0b00111100, 0b00000011, 0b11000000, 0b00000000, 
    0b01111100, 0b00000011, 0b11000000, 0b00000000, 
    0b00000000, 0b00000111, 0b11000000, 0b00000000, 
    0b00000000, 0b00001111, 0b10000000, 0b00000000, 
    0b00000001, 0b11111111, 0b10000000, 0b00000000, 
    0b00000001, 0b11111111, 0b00000000, 0b00000000, 
    0b00000001, 0b11111111, 0b00000000, 0b00000000, 
    0b00000001, 0b11111111, 0b10000000, 0b00000000, 
    0b00000000, 0b00000111, 0b11000000, 0b00000000, 
    0b00000000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111100, 0b00000111, 0b11000000, 0b00000000, 
    0b00111110, 0b00001111, 0b11000000, 0b00000000, 
    0b00111111, 0b11111111, 0b10000000, 0b00000000, 
    0b00011111, 0b11111111, 0b00000000, 0b00000000, 
    0b00001111, 0b11111110, 0b00000000, 0b00000000, 
    0b00000011, 0b11111000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter num_four={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00001110, 0b00000000, 0b00000000, 
    0b00000000, 0b00011110, 0b00000000, 0b00000000, 
    0b00000000, 0b00111110, 0b00000000, 0b00000000, 
    0b00000000, 0b01111110, 0b00000000, 0b00000000, 
    0b00000000, 0b11111110, 0b00000000, 0b00000000, 
    0b00000000, 0b11111110, 0b00000000, 0b00000000, 
    0b00000001, 0b11111110, 0b00000000, 0b00000000, 
    0b00000011, 0b11101110, 0b00000000, 0b00000000, 
    0b00000111, 0b11001110, 0b00000000, 0b00000000, 
    0b00000111, 0b10001110, 0b00000000, 0b00000000, 
    0b00001111, 0b10001110, 0b00000000, 0b00000000, 
    0b00011111, 0b00001110, 0b00000000, 0b00000000, 
    0b00111110, 0b00001110, 0b00000000, 0b00000000, 
    0b00111100, 0b00001110, 0b00000000, 0b00000000, 
    0b01111100, 0b00001110, 0b00000000, 0b00000000, 
    0b11111000, 0b00001110, 0b00000000, 0b00000000, 
    0b11111111, 0b11111111, 0b11100000, 0b00000000, 
    0b11111111, 0b11111111, 0b11100000, 0b00000000, 
    0b11111111, 0b11111111, 0b11100000, 0b00000000, 
    0b00000000, 0b00001110, 0b00000000, 0b00000000, 
    0b00000000, 0b00001110, 0b00000000, 0b00000000, 
    0b00000000, 0b00001110, 0b00000000, 0b00000000, 
    0b00000000, 0b00001110, 0b00000000, 0b00000000, 
    0b00000000, 0b00001110, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter num_five={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b10000000, 0b00000000, 
    0b00011111, 0b11111111, 0b10000000, 0b00000000, 
    0b00111111, 0b11111111, 0b10000000, 0b00000000, 
    0b00111111, 0b11111111, 0b10000000, 0b00000000, 
    0b00111100, 0b00000000, 0b00000000, 0b00000000, 
    0b00111100, 0b00000000, 0b00000000, 0b00000000, 
    0b00111100, 0b00000000, 0b00000000, 0b00000000, 
    0b00111100, 0b00000000, 0b00000000, 0b00000000, 
    0b00111101, 0b11111100, 0b00000000, 0b00000000, 
    0b00111111, 0b11111110, 0b00000000, 0b00000000, 
    0b00111111, 0b11111111, 0b00000000, 0b00000000, 
    0b00111111, 0b11111111, 0b10000000, 0b00000000, 
    0b00111110, 0b00001111, 0b11000000, 0b00000000, 
    0b01111100, 0b00000111, 0b11000000, 0b00000000, 
    0b00000000, 0b00000011, 0b11000000, 0b00000000, 
    0b00000000, 0b00000011, 0b11000000, 0b00000000, 
    0b00000000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111100, 0b00000111, 0b11000000, 0b00000000, 
    0b00111110, 0b00001111, 0b10000000, 0b00000000, 
    0b00111111, 0b11111111, 0b10000000, 0b00000000, 
    0b00011111, 0b11111111, 0b00000000, 0b00000000, 
    0b00001111, 0b11111110, 0b00000000, 0b00000000, 
    0b00000011, 0b11111000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter num_six={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11111100, 0b00000000, 0b00000000, 
    0b00000111, 0b11111111, 0b00000000, 0b00000000, 
    0b00001111, 0b11111111, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b10000000, 0b00000000, 
    0b00011111, 0b00000111, 0b10000000, 0b00000000, 
    0b00111110, 0b00000111, 0b11000000, 0b00000000, 
    0b00111100, 0b00000011, 0b11000000, 0b00000000, 
    0b01111100, 0b00000000, 0b00000000, 0b00000000, 
    0b01111000, 0b11111000, 0b00000000, 0b00000000, 
    0b01111011, 0b11111110, 0b00000000, 0b00000000, 
    0b01111111, 0b11111111, 0b00000000, 0b00000000, 
    0b01111111, 0b11111111, 0b10000000, 0b00000000, 
    0b01111111, 0b00001111, 0b11000000, 0b00000000, 
    0b01111110, 0b00000111, 0b11000000, 0b00000000, 
    0b01111100, 0b00000011, 0b11000000, 0b00000000, 
    0b01111100, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111100, 0b00000011, 0b11000000, 0b00000000, 
    0b00111100, 0b00000011, 0b11000000, 0b00000000, 
    0b00111100, 0b00000111, 0b11000000, 0b00000000, 
    0b00111111, 0b00001111, 0b10000000, 0b00000000, 
    0b00011111, 0b11111111, 0b10000000, 0b00000000, 
    0b00001111, 0b11111111, 0b00000000, 0b00000000, 
    0b00000111, 0b11111110, 0b00000000, 0b00000000, 
    0b00000001, 0b11111000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter num_seven={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b11111111, 0b11111111, 0b10000000, 0b00000000, 
    0b11111111, 0b11111111, 0b10000000, 0b00000000, 
    0b11111111, 0b11111111, 0b10000000, 0b00000000, 
    0b11111111, 0b11111111, 0b10000000, 0b00000000, 
    0b00000000, 0b00001111, 0b00000000, 0b00000000, 
    0b00000000, 0b00001111, 0b00000000, 0b00000000, 
    0b00000000, 0b00011111, 0b00000000, 0b00000000, 
    0b00000000, 0b00011110, 0b00000000, 0b00000000, 
    0b00000000, 0b00111110, 0b00000000, 0b00000000, 
    0b00000000, 0b00111100, 0b00000000, 0b00000000, 
    0b00000000, 0b00111100, 0b00000000, 0b00000000, 
    0b00000000, 0b01111100, 0b00000000, 0b00000000, 
    0b00000000, 0b01111000, 0b00000000, 0b00000000, 
    0b00000000, 0b11111000, 0b00000000, 0b00000000, 
    0b00000000, 0b11110000, 0b00000000, 0b00000000, 
    0b00000001, 0b11110000, 0b00000000, 0b00000000, 
    0b00000001, 0b11110000, 0b00000000, 0b00000000, 
    0b00000001, 0b11100000, 0b00000000, 0b00000000, 
    0b00000011, 0b11100000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000000, 0b00000000, 0b00000000, 
    0b00000111, 0b11000000, 0b00000000, 0b00000000, 
    0b00000111, 0b11000000, 0b00000000, 0b00000000, 
    0b00000111, 0b10000000, 0b00000000, 0b00000000, 
    0b00001111, 0b10000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter num_eight={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000111, 0b11111100, 0b00000000, 0b00000000, 
    0b00001111, 0b11111110, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b00000000, 0b00000000, 
    0b00111111, 0b10111111, 0b10000000, 0b00000000, 
    0b00111110, 0b00000111, 0b10000000, 0b00000000, 
    0b01111100, 0b00000111, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b00111100, 0b00000011, 0b11000000, 0b00000000, 
    0b00111100, 0b00000111, 0b11000000, 0b00000000, 
    0b00111110, 0b00001111, 0b10000000, 0b00000000, 
    0b00011111, 0b11111111, 0b10000000, 0b00000000, 
    0b00001111, 0b11111110, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b10000000, 0b00000000, 
    0b00111111, 0b11111111, 0b10000000, 0b00000000, 
    0b01111110, 0b00000111, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11100000, 0b00000000, 
    0b01111000, 0b00000011, 0b11100000, 0b00000000, 
    0b01111100, 0b00000011, 0b11000000, 0b00000000, 
    0b01111110, 0b00000111, 0b11000000, 0b00000000, 
    0b00111111, 0b11111111, 0b11000000, 0b00000000, 
    0b00111111, 0b11111111, 0b10000000, 0b00000000, 
    0b00001111, 0b11111110, 0b00000000, 0b00000000, 
    0b00000011, 0b11111000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter num_nine={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000011, 0b11111000, 0b00000000, 0b00000000, 
    0b00001111, 0b11111110, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b00000000, 0b00000000, 
    0b00111111, 0b11111111, 0b00000000, 0b00000000, 
    0b00111110, 0b00001111, 0b10000000, 0b00000000, 
    0b01111100, 0b00000111, 0b10000000, 0b00000000, 
    0b01111000, 0b00000111, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000011, 0b11000000, 0b00000000, 
    0b01111100, 0b00000111, 0b11000000, 0b00000000, 
    0b01111100, 0b00000111, 0b11000000, 0b00000000, 
    0b00111111, 0b00011111, 0b11000000, 0b00000000, 
    0b00111111, 0b11111111, 0b11000000, 0b00000000, 
    0b00011111, 0b11111111, 0b11000000, 0b00000000, 
    0b00000111, 0b11111011, 0b11000000, 0b00000000, 
    0b00000000, 0b11000011, 0b11000000, 0b00000000, 
    0b01111000, 0b00000111, 0b11000000, 0b00000000, 
    0b01111100, 0b00000111, 0b10000000, 0b00000000, 
    0b00111100, 0b00001111, 0b10000000, 0b00000000, 
    0b00111110, 0b00011111, 0b00000000, 0b00000000, 
    0b00111111, 0b11111111, 0b00000000, 0b00000000, 
    0b00011111, 0b11111110, 0b00000000, 0b00000000, 
    0b00001111, 0b11111100, 0b00000000, 0b00000000, 
    0b00000011, 0b11110000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter char_neg={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b01111111, 0b11111111, 0b11000000, 0b00000000, 
    0b01111111, 0b11111111, 0b11000000, 0b00000000, 
    0b01111111, 0b11111111, 0b11000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}

parameter char_dai={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000001, 0b11000000, 0b00011110, 0b00000000, 
    0b00000011, 0b11100000, 0b00011110, 0b00000000, 
    0b00000011, 0b11000000, 0b00011110, 0b00000000, 
    0b00000111, 0b11001111, 0b11111111, 0b11111100, 
    0b00001111, 0b10001111, 0b11111111, 0b11111100, 
    0b00011111, 0b00001111, 0b11111111, 0b11111100, 
    0b00111111, 0b00001111, 0b11111111, 0b11111100, 
    0b01111110, 0b11000000, 0b00011110, 0b00000000, 
    0b01111100, 0b11110000, 0b00011110, 0b00000000, 
    0b01111001, 0b11111111, 0b11111111, 0b11111110, 
    0b01110011, 0b11111111, 0b11111111, 0b11111110, 
    0b00000011, 0b11011111, 0b11111111, 0b11111110, 
    0b00000111, 0b11011111, 0b11111111, 0b11111110, 
    0b00001111, 0b10000000, 0b00000001, 0b11100000, 
    0b00011111, 0b10000000, 0b00000001, 0b11100000, 
    0b00111111, 0b10000000, 0b00000001, 0b11100000, 
    0b01111111, 0b10011111, 0b11111111, 0b11111110, 
    0b01111111, 0b10011111, 0b11111111, 0b11111110, 
    0b01111111, 0b10011111, 0b11111111, 0b11111110, 
    0b01110111, 0b10000011, 0b10000001, 0b11100000, 
    0b00000111, 0b10000111, 0b11000001, 0b11100000, 
    0b00000111, 0b10000111, 0b11000001, 0b11100000, 
    0b00000111, 0b10000011, 0b11100001, 0b11100000, 
    0b00000111, 0b10000001, 0b11110001, 0b11100000, 
    0b00000111, 0b10000000, 0b11110001, 0b11100000, 
    0b00000111, 0b10000000, 0b01110001, 0b11100000, 
    0b00000111, 0b10000000, 0b00000001, 0b11100000, 
    0b00000111, 0b10000000, 0b00111111, 0b11100000, 
    0b00000111, 0b10000000, 0b00111111, 0b11100000, 
    0b00000111, 0b10000000, 0b00111111, 0b11000000, 
    0b00000111, 0b00000000, 0b00000000, 0b00000000
}

parameter char_ding={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000111, 0b10000000, 0b00000000, 
    0b00000000, 0b00000111, 0b10000000, 0b00000000, 
    0b00000000, 0b00000111, 0b11000000, 0b00000000, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111100, 0b00000000, 0b00000000, 0b00111100, 
    0b00111100, 0b00000000, 0b00000000, 0b00111100, 
    0b00111101, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11000000, 
    0b00000011, 0b11111111, 0b11111111, 0b11000000, 
    0b00000000, 0b00000011, 0b11000000, 0b00000000, 
    0b00000001, 0b10000011, 0b11000000, 0b00000000, 
    0b00000001, 0b11000011, 0b11000000, 0b00000000, 
    0b00000011, 0b11000011, 0b11000000, 0b00000000, 
    0b00000011, 0b11000011, 0b11111111, 0b11110000, 
    0b00000011, 0b11000011, 0b11111111, 0b11110000, 
    0b00000111, 0b11000011, 0b11111111, 0b11110000, 
    0b00000111, 0b10000011, 0b11111111, 0b11110000, 
    0b00000111, 0b11000011, 0b11000000, 0b00000000, 
    0b00001111, 0b11100011, 0b11000000, 0b00000000, 
    0b00001111, 0b11110011, 0b11000000, 0b00000000, 
    0b00011111, 0b11111011, 0b11000000, 0b00000000, 
    0b00111110, 0b11111111, 0b11000000, 0b00000000, 
    0b01111110, 0b01111111, 0b11111100, 0b00000110, 
    0b01111100, 0b00011111, 0b11111111, 0b11111110, 
    0b01111000, 0b00000111, 0b11111111, 0b11111110, 
    0b01110000, 0b00000000, 0b01111111, 0b11111110, 
    0b00110000, 0b00000000, 0b00000000, 0b00000000
}

parameter char_mo={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000111, 0b10000001, 0b11100011, 0b11000000, 
    0b00000111, 0b10000001, 0b11100011, 0b11000000, 
    0b00000111, 0b10000001, 0b11100011, 0b11000000, 
    0b00000111, 0b10111111, 0b11111111, 0b11111110, 
    0b00000111, 0b10111111, 0b11111111, 0b11111110, 
    0b00000111, 0b10111111, 0b11111111, 0b11111110, 
    0b00111111, 0b11110001, 0b11100011, 0b11000000, 
    0b01111111, 0b11110001, 0b11100011, 0b11000000, 
    0b01111111, 0b11111111, 0b11111111, 0b11111000, 
    0b00111111, 0b11111111, 0b11111111, 0b11111000, 
    0b00000111, 0b10001111, 0b11111111, 0b11111000, 
    0b00001111, 0b10001111, 0b00000000, 0b01111000, 
    0b00001111, 0b11001111, 0b11111111, 0b11111000, 
    0b00001111, 0b11101111, 0b11111111, 0b11111000, 
    0b00011111, 0b11111111, 0b11111111, 0b11111000, 
    0b00011111, 0b11111111, 0b00000000, 0b01111000, 
    0b00111111, 0b11111111, 0b11111111, 0b11111000, 
    0b01111111, 0b11111111, 0b11111111, 0b11111000, 
    0b01111111, 0b10111111, 0b11111111, 0b11111000, 
    0b11111111, 0b10000000, 0b00011100, 0b00000000, 
    0b01110111, 0b10111111, 0b11111111, 0b11111110, 
    0b01100111, 0b10111111, 0b11111111, 0b11111110, 
    0b01100111, 0b10111111, 0b11111111, 0b11111110, 
    0b00000111, 0b10111111, 0b11111111, 0b11111110, 
    0b00000111, 0b10000001, 0b11111111, 0b10000000, 
    0b00000111, 0b10000011, 0b11110111, 0b11100000, 
    0b00000111, 0b10001111, 0b11100011, 0b11111000, 
    0b00000111, 0b10111111, 0b11000001, 0b11111110, 
    0b00000111, 0b10111111, 0b10000000, 0b11111110, 
    0b00000111, 0b10111100, 0b00000000, 0b00111110, 
    0b00000011, 0b10110000, 0b00000000, 0b00001100
}

parameter char_shi={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b01111000, 0b11000000, 
    0b00000000, 0b00000000, 0b01111011, 0b11000000, 
    0b00000000, 0b00000000, 0b01111011, 0b11100000, 
    0b00000000, 0b00000000, 0b01111001, 0b11110000, 
    0b00000000, 0b00000000, 0b01111000, 0b11110000, 
    0b00000000, 0b00000000, 0b01111000, 0b11110000, 
    0b01111111, 0b11111111, 0b11111111, 0b11111110, 
    0b01111111, 0b11111111, 0b11111111, 0b11111110, 
    0b01111111, 0b11111111, 0b11111111, 0b11111110, 
    0b00000000, 0b00000000, 0b01111000, 0b00000000, 
    0b00000000, 0b00000000, 0b01111000, 0b00000000, 
    0b00000000, 0b00000000, 0b01111000, 0b00000000, 
    0b00000000, 0b00000000, 0b00111000, 0b00000000, 
    0b00111111, 0b11111111, 0b10111100, 0b00000000, 
    0b00111111, 0b11111111, 0b10111100, 0b00000000, 
    0b00111111, 0b11111111, 0b10111100, 0b00000000, 
    0b00111111, 0b11111111, 0b10111100, 0b00000000, 
    0b00000000, 0b11100000, 0b00111100, 0b00000000, 
    0b00000000, 0b11100000, 0b00111110, 0b00000000, 
    0b00000000, 0b11100000, 0b00011110, 0b00000000, 
    0b00000000, 0b11100000, 0b00011110, 0b00000000, 
    0b00000000, 0b11100000, 0b00011110, 0b00001000, 
    0b00000000, 0b11100000, 0b11001111, 0b00011110, 
    0b00000000, 0b11111111, 0b11001111, 0b00011110, 
    0b00000111, 0b11111111, 0b11001111, 0b10011110, 
    0b01111111, 0b11111111, 0b11000111, 0b10011110, 
    0b01111111, 0b11111110, 0b00000111, 0b11111100, 
    0b00111111, 0b10000000, 0b00000011, 0b11111100, 
    0b00110000, 0b00000000, 0b00000001, 0b11111000, 
    0b00000000, 0b00000000, 0b00000001, 0b11111000, 
    0b00000000, 0b00000000, 0b00000000, 0b00100000
}
parameter char_ji={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00001100, 0b00000000, 0b00011110, 0b00000000, 
    0b00011110, 0b00000000, 0b00011110, 0b00000000, 
    0b00011111, 0b00000000, 0b00011110, 0b00000000, 
    0b00011111, 0b11000000, 0b00011110, 0b00000000, 
    0b00000111, 0b11100000, 0b00011110, 0b00000000, 
    0b00000011, 0b11100000, 0b00011110, 0b00000000, 
    0b00000001, 0b11100000, 0b00011110, 0b00000000, 
    0b00000000, 0b11000000, 0b00011110, 0b00000000, 
    0b00000000, 0b00000000, 0b00011110, 0b00000000, 
    0b00000000, 0b00000000, 0b00011110, 0b00000000, 
    0b01111111, 0b10011111, 0b11111111, 0b11111110, 
    0b01111111, 0b10011111, 0b11111111, 0b11111110, 
    0b01111111, 0b10011111, 0b11111111, 0b11111110, 
    0b00000111, 0b10000000, 0b00011110, 0b00000000, 
    0b00000111, 0b10000000, 0b00011110, 0b00000000, 
    0b00000111, 0b10000000, 0b00011110, 0b00000000, 
    0b00000111, 0b10000000, 0b00011110, 0b00000000, 
    0b00000111, 0b10000000, 0b00011110, 0b00000000, 
    0b00000111, 0b10000000, 0b00011110, 0b00000000, 
    0b00000111, 0b10000000, 0b00011110, 0b00000000, 
    0b00000111, 0b10000000, 0b00011110, 0b00000000, 
    0b00000111, 0b10011000, 0b00011110, 0b00000000, 
    0b00000111, 0b11111000, 0b00011110, 0b00000000, 
    0b00000111, 0b11111000, 0b00011110, 0b00000000, 
    0b00000111, 0b11111000, 0b00011110, 0b00000000, 
    0b00000111, 0b11110000, 0b00011110, 0b00000000, 
    0b00000111, 0b11100000, 0b00011110, 0b00000000, 
    0b00000111, 0b10000000, 0b00011110, 0b00000000, 
    0b00000111, 0b00000000, 0b00011110, 0b00000000, 
    0b00000010, 0b00000000, 0b00011110, 0b00000000, 
    0b00000000, 0b00000000, 0b00011110, 0b00000000
}
parameter char_suan={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000111, 0b10000000, 0b00111100, 0b00000000, 
    0b00000111, 0b10000000, 0b00111100, 0b00000000, 
    0b00001111, 0b11111111, 0b01111111, 0b11111110, 
    0b00001111, 0b11111111, 0b01111111, 0b11111110, 
    0b00011111, 0b11111111, 0b11111111, 0b11111110, 
    0b00111110, 0b01111001, 0b11110011, 0b11000000, 
    0b01111100, 0b01111001, 0b11110011, 0b11100000, 
    0b01111111, 0b11111111, 0b11111111, 0b11100000, 
    0b00111111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b10000000, 0b00000000, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b10000000, 0b00000000, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000000, 0b01111000, 0b00001111, 0b00000000, 
    0b01111111, 0b11111111, 0b11111111, 0b11111110, 
    0b01111111, 0b11111111, 0b11111111, 0b11111110, 
    0b01111111, 0b11111111, 0b11111111, 0b11111110, 
    0b00000001, 0b11110000, 0b00001111, 0b00000000, 
    0b00000011, 0b11110000, 0b00001111, 0b00000000, 
    0b00011111, 0b11100000, 0b00001111, 0b00000000, 
    0b00011111, 0b11000000, 0b00001111, 0b00000000, 
    0b00001111, 0b00000000, 0b00001111, 0b00000000, 
    0b00001100, 0b00000000, 0b00001110, 0b00000000
}
parameter char_xue={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000011, 0b00000111, 0b00000001, 0b11100000, 
    0b00001111, 0b00001111, 0b00000001, 0b11100000, 
    0b00001111, 0b10001111, 0b10000011, 0b11100000, 
    0b00000111, 0b11000111, 0b11000011, 0b11100000, 
    0b00000011, 0b11000011, 0b11000111, 0b11000000, 
    0b00000011, 0b11100011, 0b11000111, 0b11000000, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111000, 0b00000000, 0b00000000, 0b00011100, 
    0b00111001, 0b11111111, 0b11111111, 0b10011100, 
    0b00111001, 0b11111111, 0b11111111, 0b10011100, 
    0b00111001, 0b11111111, 0b11111111, 0b10011100, 
    0b00111001, 0b11111111, 0b11111111, 0b10011100, 
    0b00000000, 0b00000000, 0b01111111, 0b00000000, 
    0b00000000, 0b00000001, 0b11111100, 0b00000000, 
    0b00000000, 0b00000001, 0b11111000, 0b00000000, 
    0b00000000, 0b00000001, 0b11100000, 0b00000000, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00000000, 0b00000001, 0b11000000, 0b00000000, 
    0b00000000, 0b00000001, 0b11000000, 0b00000000, 
    0b00000000, 0b00000001, 0b11000000, 0b00000000, 
    0b00000000, 0b00000011, 0b11000000, 0b00000000, 
    0b00000000, 0b00111111, 0b11000000, 0b00000000, 
    0b00000000, 0b00111111, 0b11000000, 0b00000000, 
    0b00000000, 0b00111111, 0b11000000, 0b00000000, 
    0b00000000, 0b00111111, 0b00000000, 0b00000000
}
parameter char_xi={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00011111, 0b11111111, 0b11111111, 0b11110000, 
    0b00011111, 0b11111111, 0b11111111, 0b11110000, 
    0b00011111, 0b11111111, 0b11111111, 0b11110000, 
    0b00001111, 0b11111111, 0b11111111, 0b11110000, 
    0b00000000, 0b00000000, 0b00000000, 0b11110000, 
    0b00000001, 0b10000000, 0b00000000, 0b11110000, 
    0b00000011, 0b11000000, 0b00000000, 0b11110000, 
    0b00000111, 0b11100000, 0b00000000, 0b11110000, 
    0b00000011, 0b11110000, 0b00000000, 0b11110000, 
    0b00000001, 0b11111000, 0b00000000, 0b11110000, 
    0b00000000, 0b11111100, 0b00000000, 0b11110000, 
    0b00000000, 0b00111110, 0b00000000, 0b11110000, 
    0b00000000, 0b00011110, 0b00000000, 0b11110000, 
    0b00000000, 0b00001100, 0b00011000, 0b11110000, 
    0b00000000, 0b00000000, 0b01111100, 0b11110000, 
    0b00000000, 0b00000001, 0b11111100, 0b11110000, 
    0b00000000, 0b00000111, 0b11111100, 0b11110000, 
    0b00000000, 0b00011111, 0b11110000, 0b11110000, 
    0b00000000, 0b11111111, 0b11000000, 0b11110000, 
    0b00000111, 0b11111111, 0b00000000, 0b11110000, 
    0b00011111, 0b11111100, 0b00000000, 0b11110000, 
    0b00011111, 0b11100000, 0b00000000, 0b11100000, 
    0b00011111, 0b10000000, 0b00000000, 0b11100000, 
    0b00011100, 0b00000000, 0b00000001, 0b11100000, 
    0b00000000, 0b00000000, 0b00000001, 0b11100000, 
    0b00000000, 0b00000000, 0b11111111, 0b11100000, 
    0b00000000, 0b00000000, 0b11111111, 0b11000000, 
    0b00000000, 0b00000000, 0b11111111, 0b11000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}
parameter char_jing={
     0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000111, 0b10000000, 0b00000000, 
    0b00000000, 0b00000111, 0b11000000, 0b00000000, 
    0b00000000, 0b00000011, 0b11000000, 0b00000000, 
    0b00011111, 0b11111111, 0b11111111, 0b11111000, 
    0b00011111, 0b11111111, 0b11111111, 0b11111000, 
    0b00011111, 0b11111111, 0b11111111, 0b11111000, 
    0b00000000, 0b11111000, 0b00011111, 0b00000000, 
    0b00000000, 0b01111000, 0b00011110, 0b00000000, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b10000000, 0b00000001, 0b11100000, 
    0b00000111, 0b10000000, 0b00000001, 0b11100000, 
    0b00000111, 0b10000000, 0b00000001, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000011, 0b11111111, 0b11111111, 0b11101000, 
    0b00000000, 0b00111110, 0b01111000, 0b00011110, 
    0b00000000, 0b01111100, 0b01111000, 0b00011110, 
    0b00000000, 0b11111100, 0b01111000, 0b00011110, 
    0b00000111, 0b11111000, 0b01111100, 0b00111110, 
    0b01111111, 0b11110000, 0b00111111, 0b11111110, 
    0b01111111, 0b11000000, 0b00111111, 0b11111100, 
    0b01111111, 0b00000000, 0b00011111, 0b11111000, 
    0b00111000, 0b00000000, 0b00000000, 0b00000000
}

parameter char_sai={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000111, 0b10000000, 0b00000000, 
    0b00000000, 0b00000111, 0b11000000, 0b00000000, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111100, 0b00111100, 0b00111000, 0b00111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00000011, 0b11111111, 0b11111111, 0b11000000, 
    0b00000011, 0b11111111, 0b11111111, 0b11000000, 
    0b00000011, 0b11111111, 0b11111111, 0b11000000, 
    0b00000011, 0b11111111, 0b11111111, 0b11000000, 
    0b00000000, 0b00111100, 0b00111000, 0b00000000, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00000011, 0b11110000, 0b00001111, 0b11000000, 
    0b00011111, 0b11111111, 0b11111111, 0b11111000, 
    0b01111111, 0b11111111, 0b11111111, 0b11111110, 
    0b01111111, 0b11111111, 0b11111111, 0b11111110, 
    0b00111001, 0b11000011, 0b11000011, 0b10011100, 
    0b00000001, 0b11000011, 0b11000011, 0b10000000, 
    0b00000001, 0b11000011, 0b10000011, 0b10000000, 
    0b00000001, 0b11000111, 0b10000011, 0b10000000, 
    0b00000001, 0b11000111, 0b11110011, 0b10000000, 
    0b00000001, 0b11001111, 0b11111111, 0b10000000, 
    0b00000000, 0b00111111, 0b11111111, 0b11000000, 
    0b00001111, 0b11111111, 0b00111111, 0b11110000, 
    0b00011111, 0b11111100, 0b00000111, 0b11110000, 
    0b00001111, 0b11111000, 0b00000001, 0b11110000, 
    0b00001111, 0b00000000, 0b00000000, 0b01100000
}

parameter char_yan={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b01111000, 0b00000000, 
    0b00111100, 0b00000000, 0b01111000, 0b00000000, 
    0b01111110, 0b00111111, 0b11111111, 0b11111110, 
    0b00111111, 0b00111111, 0b11111111, 0b11111110, 
    0b00011111, 0b10111111, 0b11111111, 0b11111110, 
    0b00001111, 0b11111111, 0b11111111, 0b11111110, 
    0b00000111, 0b11111000, 0b00000000, 0b00011110, 
    0b00000011, 0b10111111, 0b11111111, 0b11111110, 
    0b00110000, 0b00111111, 0b11111111, 0b11111110, 
    0b01111000, 0b00111111, 0b11111111, 0b11111100, 
    0b01111110, 0b00000000, 0b00111100, 0b00000000, 
    0b01111111, 0b00011111, 0b11111111, 0b11111000, 
    0b00011111, 0b10011111, 0b11111111, 0b11111000, 
    0b00001111, 0b10011111, 0b11111111, 0b11111000, 
    0b00000111, 0b10011111, 0b11111111, 0b11111000, 
    0b00000011, 0b00011110, 0b00111100, 0b00111000, 
    0b00000000, 0b00011111, 0b11111111, 0b11111000, 
    0b00000011, 0b10011111, 0b11111111, 0b11111000, 
    0b00000011, 0b11011111, 0b11111111, 0b11111000, 
    0b00000111, 0b11011110, 0b00111100, 0b00111000, 
    0b00000111, 0b10011110, 0b00111100, 0b00111000, 
    0b00000111, 0b10011111, 0b11111111, 0b11111000, 
    0b00001111, 0b00011111, 0b11111111, 0b11111000, 
    0b00001111, 0b00011111, 0b11111111, 0b11111000, 
    0b00011110, 0b00000001, 0b11000011, 0b10000000, 
    0b00011110, 0b00000111, 0b11100011, 0b11100000, 
    0b00111100, 0b00011111, 0b11100011, 0b11111000, 
    0b00111100, 0b01111111, 0b10000001, 0b11111110, 
    0b01111100, 0b11111111, 0b00000000, 0b01111111, 
    0b00111000, 0b01111100, 0b00000000, 0b00011110, 
    0b00000000, 0b00110000, 0b00000000, 0b00000100
}
parameter char_shi2={
     0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000111, 0b11111111, 0b11111111, 0b11100000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00111111, 0b11111111, 0b11111111, 0b11111100, 
    0b00000000, 0b00000011, 0b11000000, 0b00000000, 
    0b00000000, 0b00000011, 0b11000001, 0b10000000, 
    0b00000011, 0b11000011, 0b11000111, 0b10000000, 
    0b00000011, 0b11000011, 0b11000011, 0b11000000, 
    0b00000011, 0b11000011, 0b11000011, 0b11100000, 
    0b00000111, 0b10000011, 0b11000001, 0b11100000, 
    0b00000111, 0b10000011, 0b11000001, 0b11110000, 
    0b00001111, 0b10000011, 0b11000000, 0b11110000, 
    0b00001111, 0b00000011, 0b11000000, 0b11111000, 
    0b00011111, 0b00000011, 0b11000000, 0b01111000, 
    0b00111110, 0b00000011, 0b11000000, 0b01111100, 
    0b00111110, 0b00000011, 0b11000000, 0b00111100, 
    0b01111100, 0b00000011, 0b11000000, 0b00111110, 
    0b01111000, 0b01111111, 0b11000000, 0b00011110, 
    0b00011000, 0b01111111, 0b11000000, 0b00011000, 
    0b00000000, 0b01111111, 0b10000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b00000000
}
parameter char_dui={
     0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000000, 0b00000000, 0b00000000, 0b11110000, 
    0b00000000, 0b00000000, 0b00000000, 0b11110000, 
    0b00000000, 0b00000000, 0b00000000, 0b11110000, 
    0b00111111, 0b11111100, 0b00000000, 0b11110000, 
    0b00111111, 0b11111100, 0b00000000, 0b11110000, 
    0b00111111, 0b11111100, 0b00000000, 0b11110000, 
    0b00111111, 0b11111101, 0b11111111, 0b11111110, 
    0b00000000, 0b00011101, 0b11111111, 0b11111110, 
    0b00011000, 0b00111101, 0b11111111, 0b11111110, 
    0b00111000, 0b00111101, 0b11111111, 0b11111110, 
    0b00111100, 0b00111100, 0b00000000, 0b11110000, 
    0b00111110, 0b00111100, 0b00000000, 0b11110000, 
    0b00011111, 0b00111000, 0b11000000, 0b11110000, 
    0b00001111, 0b11111001, 0b11100000, 0b11110000, 
    0b00001111, 0b11111001, 0b11100000, 0b11110000, 
    0b00000111, 0b11110001, 0b11110000, 0b11110000, 
    0b00000011, 0b11110000, 0b11111000, 0b11110000, 
    0b00000001, 0b11110000, 0b01111000, 0b11110000, 
    0b00000001, 0b11111000, 0b01111100, 0b11110000, 
    0b00000011, 0b11111000, 0b00111110, 0b11110000, 
    0b00000111, 0b11111100, 0b00011110, 0b11110000, 
    0b00000111, 0b11111110, 0b00011000, 0b11110000, 
    0b00001111, 0b10011110, 0b00000000, 0b11110000, 
    0b00011111, 0b00011110, 0b00000000, 0b11110000, 
    0b00111110, 0b00001100, 0b00000000, 0b11110000, 
    0b01111100, 0b00000000, 0b00000000, 0b11110000, 
    0b01111000, 0b00000000, 0b00000000, 0b11110000, 
    0b01110000, 0b00000000, 0b01111111, 0b11100000, 
    0b00100000, 0b00000000, 0b01111111, 0b11100000, 
    0b00000000, 0b00000000, 0b00111111, 0b11100000, 
    0b00000000, 0b00000000, 0b00111111, 0b10000000
}

parameter char_cuo={
    0b00000000, 0b00000000, 0b00000000, 0b00000000, 
    0b00000111, 0b00000000, 0b01110000, 0b11100000, 
    0b00001111, 0b00000000, 0b01110000, 0b11100000, 
    0b00001111, 0b00000000, 0b01110000, 0b11100000, 
    0b00001111, 0b00000000, 0b01110000, 0b11100000, 
    0b00011111, 0b11111111, 0b11111111, 0b11111110, 
    0b00011111, 0b11111111, 0b11111111, 0b11111110, 
    0b00011111, 0b11111111, 0b11111111, 0b11111110, 
    0b00111100, 0b00000000, 0b01110000, 0b11100000, 
    0b00111100, 0b00000000, 0b01110000, 0b11100000, 
    0b01111000, 0b00000000, 0b01110000, 0b11100000, 
    0b11111111, 0b11111111, 0b11111111, 0b11111110, 
    0b11111111, 0b11111111, 0b11111111, 0b11111110, 
    0b01111111, 0b11111111, 0b11111111, 0b11111110, 
    0b00001111, 0b11110000, 0b00000000, 0b00000000, 
    0b00000011, 0b11000001, 0b11111111, 0b11111000, 
    0b00000011, 0b11000001, 0b11111111, 0b11111000, 
    0b00111111, 0b11111101, 0b11111111, 0b11111000, 
    0b00111111, 0b11111101, 0b11111111, 0b11111000, 
    0b00111111, 0b11111101, 0b11000000, 0b00111000, 
    0b00111111, 0b11111101, 0b11000000, 0b00111000, 
    0b00000011, 0b11000001, 0b11111111, 0b11111000, 
    0b00000011, 0b11000001, 0b11111111, 0b11111000, 
    0b00000011, 0b11000001, 0b11111111, 0b11111000, 
    0b00000011, 0b11000001, 0b11000000, 0b00111000, 
    0b00000011, 0b11011101, 0b11000000, 0b00111000, 
    0b00000011, 0b11111111, 0b11000000, 0b00111000, 
    0b00000111, 0b11111111, 0b11111111, 0b11111000, 
    0b00000111, 0b11111001, 0b11111111, 0b11111000, 
    0b00000111, 0b11100001, 0b11111111, 0b11111000, 
    0b00000011, 0b00000001, 0b11000000, 0b00111000, 
    0b00000000, 0b00000001, 0b11000000, 0b00111000
}
`endif // VGA_CHAR_PARAMS_VH