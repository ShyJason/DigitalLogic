// vga_char_params.vh
`ifndef VGA_CHAR_PARAMS_VH
`define VGA_CHAR_PARAMS_VH

//num_zero- num_nine: 32x32 pixel font for numbers 0-9

//char_dai:待
//char_ding:定
//char_mo:模
//char_shi:式
//char_ji:计
//char_suan:算
//char_xue:学
//char_xi:习
//char_yan:演
//char_shi2:示
//char_dui:对
//char_cuo:错
//char_guan:关
//char_ji2:机

parameter char_none={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter num_zero={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter num_one={
     8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b01111011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b01100011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter num_two={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00011111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11100000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b10000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter num_three={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00000001, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00000001, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter num_four={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00011110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b01111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11101110, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11001110, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10001110, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b10001110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00111110, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b01111100, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b11111000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter num_five={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111101, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter num_six={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b01111011, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b01111111, 8'b00001111, 8'b11000000, 8'b00000000, 
    8'b01111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter num_seven={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b11111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00011111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00011110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b01111100, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11100000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11100000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b10000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter num_eight={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b10111111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b01111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11100000, 8'b00000000, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111110, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter num_nine={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00111110, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b01111000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b00011111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000111, 8'b11111011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b11000011, 8'b11000000, 8'b00000000, 
    8'b01111000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b01111100, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00111100, 8'b00001111, 8'b10000000, 8'b00000000, 
    8'b00111110, 8'b00011111, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter char_neg={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter char_A={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11011110, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11011111, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11011111, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10001111, 8'b00000000, 8'b00000000, 
    8'b00001111, 8'b10001111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00001111, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00011111, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00011110, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b01111100, 8'b00000001, 8'b11110000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b11110000, 8'b00000000, 
    8'b11111000, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b11111000, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b11110000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b11110000, 8'b00000000, 8'b01111100, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter char_B={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000001, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000001, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000001, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11111000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter char_C={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00000011, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11111000, 8'b00000000, 
    8'b00011111, 8'b10000001, 8'b11111000, 8'b00000000, 
    8'b00111111, 8'b00000000, 8'b01111100, 8'b00000000, 
    8'b00111110, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b01111000, 8'b00000000, 8'b00011100, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00111110, 8'b00000000, 
    8'b01111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111110, 8'b00000000, 8'b01111100, 8'b00000000, 
    8'b00111111, 8'b00000000, 8'b11111100, 8'b00000000, 
    8'b00011111, 8'b10000001, 8'b11111000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00000011, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b11111110, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter char_D={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111100, 8'b00000111, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000001, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111100, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b11111000, 8'b00000000, 
    8'b00111100, 8'b00000011, 8'b11110000, 8'b00000000, 
    8'b00111100, 8'b00001111, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter char_E={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11100000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11110000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter char_F={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter char_guan={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b01100000, 8'b00000111, 8'b10000000, 
    8'b00000001, 8'b11100000, 8'b00000111, 8'b10000000, 
    8'b00000001, 8'b11110000, 8'b00001111, 8'b00000000, 
    8'b00000000, 8'b11111000, 8'b00001111, 8'b00000000, 
    8'b00000000, 8'b01111000, 8'b00011111, 8'b00000000, 
    8'b00000000, 8'b01111100, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b00111100, 8'b00111110, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000000, 8'b00001111, 8'b11100000, 8'b00000000, 
    8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 
    8'b00000000, 8'b00011111, 8'b11111000, 8'b00000000, 
    8'b00000000, 8'b00011110, 8'b01111100, 8'b00000000, 
    8'b00000000, 8'b00111110, 8'b01111110, 8'b00000000, 
    8'b00000000, 8'b01111100, 8'b00111111, 8'b00000000, 
    8'b00000001, 8'b11111100, 8'b00011111, 8'b10000000, 
    8'b00000111, 8'b11110000, 8'b00001111, 8'b11100000, 
    8'b00011111, 8'b11100000, 8'b00000111, 8'b11111100, 
    8'b01111111, 8'b11000000, 8'b00000001, 8'b11111110, 
    8'b01111111, 8'b00000000, 8'b00000000, 8'b11111110, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00001100
}

parameter char_ji2={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11000011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b00000111, 8'b11000011, 8'b11000011, 8'b11000000, 
    8'b00000111, 8'b11100011, 8'b11000011, 8'b11000000, 
    8'b00001111, 8'b11110011, 8'b11000011, 8'b11000000, 
    8'b00001111, 8'b11111011, 8'b11000011, 8'b11000000, 
    8'b00001111, 8'b11111011, 8'b11000011, 8'b11000000, 
    8'b00011111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b00111111, 8'b11111111, 8'b11000011, 8'b11000000, 
    8'b00111111, 8'b11011011, 8'b11000011, 8'b11000000, 
    8'b01111011, 8'b11011011, 8'b11000011, 8'b11000000, 
    8'b01111011, 8'b11000011, 8'b11000011, 8'b11000000, 
    8'b01110011, 8'b11000011, 8'b11000011, 8'b11001110, 
    8'b01110011, 8'b11000011, 8'b10000011, 8'b11001110, 
    8'b01100011, 8'b11000111, 8'b10000011, 8'b11001110, 
    8'b00000011, 8'b11000111, 8'b10000011, 8'b11001110, 
    8'b00000011, 8'b11000111, 8'b10000011, 8'b11001110, 
    8'b00000011, 8'b11001111, 8'b00000011, 8'b11001110, 
    8'b00000011, 8'b11011111, 8'b00000011, 8'b11111110, 
    8'b00000011, 8'b11011111, 8'b00000011, 8'b11111110, 
    8'b00000011, 8'b11011110, 8'b00000001, 8'b11111110, 
    8'b00000011, 8'b11011110, 8'b00000000, 8'b11111100, 
    8'b00000011, 8'b10001100, 8'b00000000, 8'b00000000
}

parameter char_dai={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000001, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b00000011, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000011, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11001111, 8'b11111111, 8'b11111100, 
    8'b00001111, 8'b10001111, 8'b11111111, 8'b11111100, 
    8'b00011111, 8'b00001111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b00001111, 8'b11111111, 8'b11111100, 
    8'b01111110, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b01111100, 8'b11110000, 8'b00011110, 8'b00000000, 
    8'b01111001, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01110011, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00000011, 8'b11011111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b11011111, 8'b11111111, 8'b11111110, 
    8'b00001111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00011111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00111111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01110111, 8'b10000011, 8'b10000001, 8'b11100000, 
    8'b00000111, 8'b10000111, 8'b11000001, 8'b11100000, 
    8'b00000111, 8'b10000111, 8'b11000001, 8'b11100000, 
    8'b00000111, 8'b10000011, 8'b11100001, 8'b11100000, 
    8'b00000111, 8'b10000001, 8'b11110001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b11110001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b01110001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00111111, 8'b11000000, 
    8'b00000111, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter char_ding={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 
    8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 
    8'b00111101, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000001, 8'b10000011, 8'b11000000, 8'b00000000, 
    8'b00000001, 8'b11000011, 8'b11000000, 8'b00000000, 
    8'b00000011, 8'b11000011, 8'b11000000, 8'b00000000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11110000, 
    8'b00000011, 8'b11000011, 8'b11111111, 8'b11110000, 
    8'b00000111, 8'b11000011, 8'b11111111, 8'b11110000, 
    8'b00000111, 8'b10000011, 8'b11111111, 8'b11110000, 
    8'b00000111, 8'b11000011, 8'b11000000, 8'b00000000, 
    8'b00001111, 8'b11100011, 8'b11000000, 8'b00000000, 
    8'b00001111, 8'b11110011, 8'b11000000, 8'b00000000, 
    8'b00011111, 8'b11111011, 8'b11000000, 8'b00000000, 
    8'b00111110, 8'b11111111, 8'b11000000, 8'b00000000, 
    8'b01111110, 8'b01111111, 8'b11111100, 8'b00000110, 
    8'b01111100, 8'b00011111, 8'b11111111, 8'b11111110, 
    8'b01111000, 8'b00000111, 8'b11111111, 8'b11111110, 
    8'b01110000, 8'b00000000, 8'b01111111, 8'b11111110, 
    8'b00110000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter char_mo={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10000001, 8'b11100011, 8'b11000000, 
    8'b00000111, 8'b10000001, 8'b11100011, 8'b11000000, 
    8'b00000111, 8'b10000001, 8'b11100011, 8'b11000000, 
    8'b00000111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00111111, 8'b11110001, 8'b11100011, 8'b11000000, 
    8'b01111111, 8'b11110001, 8'b11100011, 8'b11000000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b10001111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b10001111, 8'b00000000, 8'b01111000, 
    8'b00001111, 8'b11001111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b11101111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b00000000, 8'b01111000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b01111111, 8'b10111111, 8'b11111111, 8'b11111000, 
    8'b11111111, 8'b10000000, 8'b00011100, 8'b00000000, 
    8'b01110111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b01100111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b01100111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10000001, 8'b11111111, 8'b10000000, 
    8'b00000111, 8'b10000011, 8'b11110111, 8'b11100000, 
    8'b00000111, 8'b10001111, 8'b11100011, 8'b11111000, 
    8'b00000111, 8'b10111111, 8'b11000001, 8'b11111110, 
    8'b00000111, 8'b10111111, 8'b10000000, 8'b11111110, 
    8'b00000111, 8'b10111100, 8'b00000000, 8'b00111110, 
    8'b00000011, 8'b10110000, 8'b00000000, 8'b00001100
}

parameter char_shi={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b11000000, 
    8'b00000000, 8'b00000000, 8'b01111011, 8'b11000000, 
    8'b00000000, 8'b00000000, 8'b01111011, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b01111001, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b11110000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00111000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10111100, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10111100, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10111100, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b10111100, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00111100, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00111110, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b11100000, 8'b00011110, 8'b00001000, 
    8'b00000000, 8'b11100000, 8'b11001111, 8'b00011110, 
    8'b00000000, 8'b11111111, 8'b11001111, 8'b00011110, 
    8'b00000111, 8'b11111111, 8'b11001111, 8'b10011110, 
    8'b01111111, 8'b11111111, 8'b11000111, 8'b10011110, 
    8'b01111111, 8'b11111110, 8'b00000111, 8'b11111100, 
    8'b00111111, 8'b10000000, 8'b00000011, 8'b11111100, 
    8'b00110000, 8'b00000000, 8'b00000001, 8'b11111000, 
    8'b00000000, 8'b00000000, 8'b00000001, 8'b11111000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00100000
}
parameter char_ji={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00001100, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00011110, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00011111, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00011111, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000011, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000001, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b11000000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b10011111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10011000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11111000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11111000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11111000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11110000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b11100000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00011110, 8'b00000000, 
    8'b00000111, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00000010, 8'b00000000, 8'b00011110, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00011110, 8'b00000000
}
parameter char_suan={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00111100, 8'b00000000, 
    8'b00000111, 8'b10000000, 8'b00111100, 8'b00000000, 
    8'b00001111, 8'b11111111, 8'b01111111, 8'b11111110, 
    8'b00001111, 8'b11111111, 8'b01111111, 8'b11111110, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00111110, 8'b01111001, 8'b11110011, 8'b11000000, 
    8'b01111100, 8'b01111001, 8'b11110011, 8'b11100000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000000, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000000, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000000, 8'b01111000, 8'b00001111, 8'b00000000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00000001, 8'b11110000, 8'b00001111, 8'b00000000, 
    8'b00000011, 8'b11110000, 8'b00001111, 8'b00000000, 
    8'b00011111, 8'b11100000, 8'b00001111, 8'b00000000, 
    8'b00011111, 8'b11000000, 8'b00001111, 8'b00000000, 
    8'b00001111, 8'b00000000, 8'b00001111, 8'b00000000, 
    8'b00001100, 8'b00000000, 8'b00001110, 8'b00000000
}
parameter char_xue={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b00000111, 8'b00000001, 8'b11100000, 
    8'b00001111, 8'b00001111, 8'b00000001, 8'b11100000, 
    8'b00001111, 8'b10001111, 8'b10000011, 8'b11100000, 
    8'b00000111, 8'b11000111, 8'b11000011, 8'b11100000, 
    8'b00000011, 8'b11000011, 8'b11000111, 8'b11000000, 
    8'b00000011, 8'b11100011, 8'b11000111, 8'b11000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111000, 8'b00000000, 8'b00000000, 8'b00011100, 
    8'b00111001, 8'b11111111, 8'b11111111, 8'b10011100, 
    8'b00111001, 8'b11111111, 8'b11111111, 8'b10011100, 
    8'b00111001, 8'b11111111, 8'b11111111, 8'b10011100, 
    8'b00111001, 8'b11111111, 8'b11111111, 8'b10011100, 
    8'b00000000, 8'b00000000, 8'b01111111, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11111100, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11111000, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11100000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000000, 8'b00000001, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000001, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00111111, 8'b00000000, 8'b00000000
}
parameter char_xi={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11110000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11110000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11110000, 
    8'b00001111, 8'b11111111, 8'b11111111, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b00000001, 8'b10000000, 8'b00000000, 8'b11110000, 
    8'b00000011, 8'b11000000, 8'b00000000, 8'b11110000, 
    8'b00000111, 8'b11100000, 8'b00000000, 8'b11110000, 
    8'b00000011, 8'b11110000, 8'b00000000, 8'b11110000, 
    8'b00000001, 8'b11111000, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00111110, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00011110, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00001100, 8'b00011000, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b01111100, 8'b11110000, 
    8'b00000000, 8'b00000001, 8'b11111100, 8'b11110000, 
    8'b00000000, 8'b00000111, 8'b11111100, 8'b11110000, 
    8'b00000000, 8'b00011111, 8'b11110000, 8'b11110000, 
    8'b00000000, 8'b11111111, 8'b11000000, 8'b11110000, 
    8'b00000111, 8'b11111111, 8'b00000000, 8'b11110000, 
    8'b00011111, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00011111, 8'b11100000, 8'b00000000, 8'b11100000, 
    8'b00011111, 8'b10000000, 8'b00000000, 8'b11100000, 
    8'b00011100, 8'b00000000, 8'b00000001, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b00000001, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b11111111, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b11111111, 8'b11000000, 
    8'b00000000, 8'b00000000, 8'b11111111, 8'b11000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter char_jing={
     8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00000000, 8'b11111000, 8'b00011111, 8'b00000000, 
    8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00000111, 8'b10000000, 8'b00000001, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11101000, 
    8'b00000000, 8'b00111110, 8'b01111000, 8'b00011110, 
    8'b00000000, 8'b01111100, 8'b01111000, 8'b00011110, 
    8'b00000000, 8'b11111100, 8'b01111000, 8'b00011110, 
    8'b00000111, 8'b11111000, 8'b01111100, 8'b00111110, 
    8'b01111111, 8'b11110000, 8'b00111111, 8'b11111110, 
    8'b01111111, 8'b11000000, 8'b00111111, 8'b11111100, 
    8'b01111111, 8'b00000000, 8'b00011111, 8'b11111000, 
    8'b00111000, 8'b00000000, 8'b00000000, 8'b00000000
}

parameter char_sai={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111100, 8'b00111100, 8'b00111000, 8'b00111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000011, 8'b11111111, 8'b11111111, 8'b11000000, 
    8'b00000000, 8'b00111100, 8'b00111000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000011, 8'b11110000, 8'b00001111, 8'b11000000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00111001, 8'b11000011, 8'b11000011, 8'b10011100, 
    8'b00000001, 8'b11000011, 8'b11000011, 8'b10000000, 
    8'b00000001, 8'b11000011, 8'b10000011, 8'b10000000, 
    8'b00000001, 8'b11000111, 8'b10000011, 8'b10000000, 
    8'b00000001, 8'b11000111, 8'b11110011, 8'b10000000, 
    8'b00000001, 8'b11001111, 8'b11111111, 8'b10000000, 
    8'b00000000, 8'b00111111, 8'b11111111, 8'b11000000, 
    8'b00001111, 8'b11111111, 8'b00111111, 8'b11110000, 
    8'b00011111, 8'b11111100, 8'b00000111, 8'b11110000, 
    8'b00001111, 8'b11111000, 8'b00000001, 8'b11110000, 
    8'b00001111, 8'b00000000, 8'b00000000, 8'b01100000
}

parameter char_yan={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b00111100, 8'b00000000, 8'b01111000, 8'b00000000, 
    8'b01111110, 8'b00111111, 8'b11111111, 8'b11111110, 
    8'b00111111, 8'b00111111, 8'b11111111, 8'b11111110, 
    8'b00011111, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00001111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00000111, 8'b11111000, 8'b00000000, 8'b00011110, 
    8'b00000011, 8'b10111111, 8'b11111111, 8'b11111110, 
    8'b00110000, 8'b00111111, 8'b11111111, 8'b11111110, 
    8'b01111000, 8'b00111111, 8'b11111111, 8'b11111100, 
    8'b01111110, 8'b00000000, 8'b00111100, 8'b00000000, 
    8'b01111111, 8'b00011111, 8'b11111111, 8'b11111000, 
    8'b00011111, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b00011110, 8'b00111100, 8'b00111000, 
    8'b00000000, 8'b00011111, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11011111, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b11011110, 8'b00111100, 8'b00111000, 
    8'b00000111, 8'b10011110, 8'b00111100, 8'b00111000, 
    8'b00000111, 8'b10011111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b00011111, 8'b11111111, 8'b11111000, 
    8'b00001111, 8'b00011111, 8'b11111111, 8'b11111000, 
    8'b00011110, 8'b00000001, 8'b11000011, 8'b10000000, 
    8'b00011110, 8'b00000111, 8'b11100011, 8'b11100000, 
    8'b00111100, 8'b00011111, 8'b11100011, 8'b11111000, 
    8'b00111100, 8'b01111111, 8'b10000001, 8'b11111110, 
    8'b01111100, 8'b11111111, 8'b00000000, 8'b01111111, 
    8'b00111000, 8'b01111100, 8'b00000000, 8'b00011110, 
    8'b00000000, 8'b00110000, 8'b00000000, 8'b00000100
}
parameter char_shi2={
     8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00111111, 8'b11111111, 8'b11111111, 8'b11111100, 
    8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 
    8'b00000000, 8'b00000011, 8'b11000001, 8'b10000000, 
    8'b00000011, 8'b11000011, 8'b11000111, 8'b10000000, 
    8'b00000011, 8'b11000011, 8'b11000011, 8'b11000000, 
    8'b00000011, 8'b11000011, 8'b11000011, 8'b11100000, 
    8'b00000111, 8'b10000011, 8'b11000001, 8'b11100000, 
    8'b00000111, 8'b10000011, 8'b11000001, 8'b11110000, 
    8'b00001111, 8'b10000011, 8'b11000000, 8'b11110000, 
    8'b00001111, 8'b00000011, 8'b11000000, 8'b11111000, 
    8'b00011111, 8'b00000011, 8'b11000000, 8'b01111000, 
    8'b00111110, 8'b00000011, 8'b11000000, 8'b01111100, 
    8'b00111110, 8'b00000011, 8'b11000000, 8'b00111100, 
    8'b01111100, 8'b00000011, 8'b11000000, 8'b00111110, 
    8'b01111000, 8'b01111111, 8'b11000000, 8'b00011110, 
    8'b00011000, 8'b01111111, 8'b11000000, 8'b00011000, 
    8'b00000000, 8'b01111111, 8'b10000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000
}
parameter char_dui={
     8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b00000000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b00111111, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00111111, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00111111, 8'b11111100, 8'b00000000, 8'b11110000, 
    8'b00111111, 8'b11111101, 8'b11111111, 8'b11111110, 
    8'b00000000, 8'b00011101, 8'b11111111, 8'b11111110, 
    8'b00011000, 8'b00111101, 8'b11111111, 8'b11111110, 
    8'b00111000, 8'b00111101, 8'b11111111, 8'b11111110, 
    8'b00111100, 8'b00111100, 8'b00000000, 8'b11110000, 
    8'b00111110, 8'b00111100, 8'b00000000, 8'b11110000, 
    8'b00011111, 8'b00111000, 8'b11000000, 8'b11110000, 
    8'b00001111, 8'b11111001, 8'b11100000, 8'b11110000, 
    8'b00001111, 8'b11111001, 8'b11100000, 8'b11110000, 
    8'b00000111, 8'b11110001, 8'b11110000, 8'b11110000, 
    8'b00000011, 8'b11110000, 8'b11111000, 8'b11110000, 
    8'b00000001, 8'b11110000, 8'b01111000, 8'b11110000, 
    8'b00000001, 8'b11111000, 8'b01111100, 8'b11110000, 
    8'b00000011, 8'b11111000, 8'b00111110, 8'b11110000, 
    8'b00000111, 8'b11111100, 8'b00011110, 8'b11110000, 
    8'b00000111, 8'b11111110, 8'b00011000, 8'b11110000, 
    8'b00001111, 8'b10011110, 8'b00000000, 8'b11110000, 
    8'b00011111, 8'b00011110, 8'b00000000, 8'b11110000, 
    8'b00111110, 8'b00001100, 8'b00000000, 8'b11110000, 
    8'b01111100, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b01111000, 8'b00000000, 8'b00000000, 8'b11110000, 
    8'b01110000, 8'b00000000, 8'b01111111, 8'b11100000, 
    8'b00100000, 8'b00000000, 8'b01111111, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b00111111, 8'b11100000, 
    8'b00000000, 8'b00000000, 8'b00111111, 8'b10000000
}

parameter char_cuo={
    8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 
    8'b00000111, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00001111, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00001111, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00001111, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00011111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00111100, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b00111100, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b01111000, 8'b00000000, 8'b01110000, 8'b11100000, 
    8'b11111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b11111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b01111111, 8'b11111111, 8'b11111111, 8'b11111110, 
    8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00111111, 8'b11111101, 8'b11111111, 8'b11111000, 
    8'b00111111, 8'b11111101, 8'b11111111, 8'b11111000, 
    8'b00111111, 8'b11111101, 8'b11000000, 8'b00111000, 
    8'b00111111, 8'b11111101, 8'b11000000, 8'b00111000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11000001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b11000001, 8'b11000000, 8'b00111000, 
    8'b00000011, 8'b11011101, 8'b11000000, 8'b00111000, 
    8'b00000011, 8'b11111111, 8'b11000000, 8'b00111000, 
    8'b00000111, 8'b11111111, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b11111001, 8'b11111111, 8'b11111000, 
    8'b00000111, 8'b11100001, 8'b11111111, 8'b11111000, 
    8'b00000011, 8'b00000001, 8'b11000000, 8'b00111000, 
    8'b00000000, 8'b00000001, 8'b11000000, 8'b00111000
}
`endif // VGA_CHAR_PARAMS_VH